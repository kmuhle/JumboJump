package sprite_package is
 type sprite_block is array(0 to 15, 0 to 15) of integer range 0 to 3;

constant acorn_head_1: sprite_block :=
((0,0,0,3,3,3,3,3,3,0,0,0,0,0,1,0), 
(0,0,3,3,3,3,3,3,3,3,3,0,1,1,1,0), 
(0,0,3,3,3,3,3,3,3,3,3,3,3,1,0,0),
(0,0,0,2,2,3,3,3,3,3,3,3,3,3,0,0),
(0,0,2,2,2,3,3,3,3,3,3,3,3,3,0,0), 
(0,0,2,2,2,2,3,3,3,3,3,3,3,3,3,0), 
(0,2,2,1,1,2,2,3,3,3,3,3,3,3,3,0), 
(0,2,2,1,1,2,2,3,3,3,3,3,3,3,3,3),
(2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3), 
(2,2,2,2,1,1,2,2,2,2,3,3,3,3,3,3),
(2,1,2,2,1,2,2,1,1,2,2,3,3,3,3,3), 
(2,2,1,2,2,2,2,1,1,2,2,2,2,3,3,3), 
(2,2,2,1,2,2,2,2,2,2,2,2,2,3,3,3),
(2,2,2,2,1,2,2,2,2,2,2,2,0,3,3,0),
(2,2,2,2,2,2,2,2,2,2,0,0,0,0,0,0), 
(2,2,2,2,2,2,2,2,0,0,0,0,0,0,0,0));

constant letter_H: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,2,2,2,2,0,2,2,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,0,2,2,2,2,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant letter_i: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,2,2,2,2,0,0,0,0,0,0,0,0,0,0),
(0,0,2,1,1,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,2,2,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,1,1,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,1,1,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,1,1,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,1,1,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,1,1,2,2,0,0,0,0,0,0,0,0,0),
(0,0,2,2,2,2,2,0,0,0,0,0,0,0,0,0),
(0,0,0,2,2,2,2,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_0: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,2,2,2,2,2,0,0,0,0,0,0),
(0,0,0,0,2,2,1,1,1,2,2,0,0,0,0,0),
(0,0,0,2,2,1,1,2,2,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,1,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,1,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,1,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,2,2,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,1,1,1,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,2,2,2,2,2,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_1: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0),
(0,0,0,0,0,2,2,1,1,2,2,0,0,0,0,0),
(0,0,0,0,0,2,1,1,1,2,2,0,0,0,0,0),
(0,0,0,0,0,2,2,1,1,2,2,0,0,0,0,0),
(0,0,0,0,0,0,2,1,1,2,2,0,0,0,0,0),
(0,0,0,0,0,0,2,1,1,2,2,0,0,0,0,0),
(0,0,0,0,2,2,2,1,1,2,2,2,0,0,0,0),
(0,0,0,0,2,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_2: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,0,0,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,1,1,1,2,2,2,2,0,0,0),
(0,0,0,2,2,1,1,2,2,2,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_3: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,0,0,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,2,1,1,2,2,0,0,0),
(0,0,0,0,2,2,1,1,1,1,2,2,2,0,0,0),
(0,0,0,2,2,2,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_4: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,2,2,2,2,2,0,0,0,0,0),
(0,0,0,0,0,2,2,1,1,1,2,2,0,0,0,0),
(0,0,0,0,2,2,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,2,1,1,2,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,1,1,2,2,2,0,0,0),
(0,0,0,0,0,0,0,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_5: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,2,2,2,2,2,2,2,2,0,0,0,0,0),
(0,0,0,2,1,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,1,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,2,1,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,2,2,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant num_6: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,0,0,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,2,2,2,2,0,0,0),
(0,0,0,2,1,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_7: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,2,2,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,1,1,2,2,2,2,0,0,0),
(0,0,0,0,0,2,1,1,2,2,2,2,0,0,0,0),
(0,0,0,0,0,2,1,1,2,2,2,0,0,0,0,0),
(0,0,0,0,0,2,1,1,2,2,0,0,0,0,0,0),
(0,0,0,0,0,2,2,2,2,2,0,0,0,0,0,0),
(0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_8: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,0,0,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant num_9: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,0,0,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,0,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,1,1,1,1,1,2,2,0,0,0),
(0,0,0,2,2,2,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,1,1,2,2,2,1,1,2,2,0,0,0),
(0,0,0,2,2,1,1,1,1,1,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0),
(0,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant jumbo_box_1: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2), 
(0,0,0,0,0,0,0,1,1,1,1,1,0,0,2,2), 
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,2,2), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,2,2), 
(2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2), 
(2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2), 
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant jumbo_box_2: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,2,2,2,2,2,0,0,0,0,0,0,0,0,0), 
(0,2,2,2,2,2,2,1,1,1,1,0,0,0,0,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,0,0,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,1,0,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,0),
(2,2,2,2,2,2,2,2,1,1,3,3,1,1,1,0),
(2,2,2,2,2,2,2,1,1,1,3,3,1,1,1,1),
(2,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1),
(2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1),
(2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1),
(2,2,2,2,1,1,1,1,1,1,3,1,1,1,1,1));

constant jumbo_box_3: sprite_block :=
((0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,0,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,2,1,2,1,2,0,0,0,0,0,0,0,0));

constant jumbo_box_4: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,3,3,0,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,0,0,0,1,1,1,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,2,1,2,1,2,0,0,0,0,0,0,0,0));

constant jumbo_box_2_dead: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,2,2,2,2,2,0,0,0,0,0,0,0,0,0), 
(0,2,2,2,2,2,2,1,1,1,1,0,0,0,0,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,0,0,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,1,0,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,0), 
(2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,0),
(2,2,2,2,2,2,2,2,1,1,3,3,3,1,1,0),
(2,2,2,2,2,2,2,1,1,1,3,1,3,1,1,1),
(2,2,2,2,2,2,2,1,1,1,3,3,3,1,1,1),
(2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1),
(2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1),
(2,2,2,2,1,1,1,1,3,3,3,3,1,1,1,1));

constant jumbo_box_4_dead: sprite_block :=
((1,1,1,1,1,1,1,1,3,1,1,3,3,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,3,0,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,0,0,0,1,1,1,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,2,1,2,1,2,0,0,0,0,0,0,0,0));


constant jumbo_walk_1_box_3: sprite_block :=
((0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,0,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,1,2,1,2,1,2,0,0,0,0,0,0,0));


constant jumbo_walk_1_box_4: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,3,3,0,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,0,0,0,1,1,1,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,1,2,1,2,1,2,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant jumbo_walk_2_box_3: sprite_block :=
((0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,0,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,2,1,2,1,2,0,0,0,0,0,0,0,0,0));


constant jumbo_walk_2_box_4: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,3,3,0,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,0,0,0,1,1,1,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,2,1,2,1,2,0,0,0,0,0,0,0,0,0,0));

constant cloud_left: sprite_block:=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,2,2,2,2,2),
(0,0,0,0,0,0,0,0,0,1,2,2,2,2,2,2),
(0,0,0,0,0,0,0,0,1,2,2,2,2,2,2,2),
(0,0,0,0,0,0,0,0,1,2,2,2,2,2,2,2),
(0,0,0,0,0,0,1,1,1,2,2,2,2,2,2,2),
(0,0,0,0,0,1,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,0,1,2,2,2,2,2,2,2,2,2,2),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1));

constant cloud_right: sprite_block:=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(2,2,2,2,2,2,1,1,0,0,0,0,0,0,0,0),
(2,2,2,2,2,2,2,1,0,0,0,0,0,0,0,0),
(2,2,2,2,2,2,2,1,1,1,0,0,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0),
(2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0));


constant ground_2: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant brown_c2_r6: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,1,1,1,0,0,1,1,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,1));


constant brown_c2_r7: sprite_block :=
((0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,1),
(0,0,0,0,0,0,0,0,1,1,1,1,0,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));




constant brown_c3_r2: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant brown_c3_r3: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1));


constant brown_c3_r4: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1));

constant brown_c3_r5: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1),
(0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1),
(0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,1,1,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant brown_c3_r6: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,1,1,1,0,1,1,0,0,0),
(0,0,0,0,0,0,0,1,1,0,0,0,1,1,1,0),
(1,0,0,0,0,0,0,1,1,0,0,0,0,1,1,0),
(1,0,0,0,0,0,0,0,1,0,0,0,0,0,1,1),
(1,0,0,0,0,0,0,0,1,0,0,0,0,0,1,1));

constant brown_c3_r7: sprite_block :=
((0,0,0,0,0,0,0,0,1,0,0,0,0,1,1,0),
(0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0),
(1,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,0,0,1,0,0,1,1,1,0,0),
(1,1,0,0,0,0,0,0,1,0,0,0,1,1,0,0),
(1,1,0,0,0,0,0,0,1,0,0,0,0,1,1,0),
(1,1,0,0,0,0,0,0,1,0,0,0,0,1,1,1),
(1,0,0,0,0,0,0,1,1,0,0,0,0,0,1,1),
(0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant brown_c4_r1 : sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1),
(0,0,0,0,0,0,1,0,0,1,0,1,1,1,1,0),
(0,0,0,0,1,1,1,1,1,1,0,1,0,0,0,0),
(0,0,0,1,0,0,1,1,0,0,0,0,0,0,0,0));

constant brown_c4_r2: sprite_block :=
((0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,1,1,0,1,0,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1),
(0,1,0,0,0,0,0,0,0,1,1,1,1,0,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,0,0,1,0),
(0,0,0,0,1,1,0,0,0,1,0,0,1,0,1,0),
(0,0,0,0,1,1,0,0,0,0,1,0,1,1,1,0),
(0,0,0,1,1,0,1,1,0,0,1,0,0,1,1,1),
(1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,0),
(0,0,0,0,0,1,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,1,1,0,0,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,1,1,0,0,1,1,1,0),
(1,1,1,1,1,0,0,0,1,0,0,0,0,1,0,0),
(0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1));


constant brown_c4_r3: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1),
(0,1,1,1,1,1,1,1,1,0,0,1,0,0,0,1),
(0,0,1,1,1,1,1,1,1,1,0,0,1,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,0,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1));

constant brown_c4_r4: sprite_block :=
((0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,1,0,0,0,1,1,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant brown_c4_r5: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,0,0,0,0,1,1,1,1),
(0,0,0,1,1,0,0,0,1,0,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(0,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1),
(0,0,0,1,1,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1));

constant brown_c4_r6: sprite_block :=
((0,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,1,1,1,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,1,1,1,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,1,1,1,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant brown_c4_r7: sprite_block :=
((0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,1),
(0,0,0,0,0,0,0,1,1,0,0,0,0,0,1,1),
(1,0,0,0,0,0,0,0,1,1,1,0,0,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant brown_c5_r1: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,0,1,1,1,0,1,0,0,0,0,0,0,0,0,0),
(0,1,0,0,0,1,0,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,1,0,1,1,0,1,0,0,0,0));


constant brown_c5_r2: sprite_block :=
((0,0,0,0,0,0,0,0,0,1,1,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,1,1,1,0,0,0,0,0,0,0,0,1,1,1),
(1,1,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,0,1,0,1,1,0,1,1,0,0,0,0,0,0),
(0,1,1,0,0,1,0,0,0,1,1,0,0,0,0,0),
(0,1,1,0,0,1,0,1,1,0,1,1,0,0,0,1),
(0,0,1,1,1,1,1,0,0,0,1,0,0,1,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,0,0,0,1,0,0,0,0,0,0,0,0),
(0,0,1,0,0,0,0,1,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0));

constant brown_c5_r3: sprite_block :=
((1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1),
(1,1,1,1,1,1,1,1,0,0,1,0,0,0,1,1),
(1,1,1,1,1,1,1,1,1,0,1,1,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0));


constant brown_c5_r4: sprite_block :=
((1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
--(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant brown_c5_r5: sprite_block :=
((1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,1,1,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1),
(1,1,1,1,0,0,0,0,0,0,0,0,1,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1));

constant brown_c5_r6: sprite_block :=
((1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0),
(1,1,1,1,0,0,0,0,0,0,0,1,1,1,0,0),
(1,1,1,1,0,0,0,0,0,1,1,1,0,0,0,0),
(1,1,1,1,0,0,0,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant brown_c5_r7: sprite_block :=
((1,1,0,0,0,0,0,1,1,0,0,0,1,0,1,1),
(1,1,0,0,0,0,0,1,1,0,0,0,1,0,0,1),
(1,1,0,0,0,0,0,0,1,0,0,0,0,0,0,1),
(1,1,0,0,0,0,0,0,1,1,0,1,0,0,0,1),
(1,1,0,0,0,0,0,0,1,1,0,1,0,0,0,0),
(1,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant brown_c6_r2: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant brown_c6_r3: sprite_block :=
((1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0));

constant brown_c6_r4: sprite_block :=
((1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0));

constant brown_c6_r5: sprite_block :=
((0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant brown_c6_r6: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,0,0,0,0,1,1,0,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,1,1,0,0),
(0,0,0,0,0,1,0,0,0,0,0,0,1,1,1,0),
(0,0,0,0,1,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,1));

constant brown_c6_r7: sprite_block :=
((0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,1),
(1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0),
(1,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0),
(1,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0),
(1,1,1,0,0,0,0,0,0,0,0,0,1,0,0,0),
(1,1,1,0,0,0,0,0,0,0,0,0,1,0,0,0),
(0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0),
(0,1,0,0,0,0,0,0,0,0,0,1,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant brown_c7_r6: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0));

constant brown_c7_r7: sprite_block :=
((1,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
(0,1,1,0,0,0,1,0,0,0,0,0,0,0,0,0),
(0,0,1,1,0,0,1,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,0,1,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant s_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1));

constant s_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0));


constant s_bottom_left: sprite_block :=
((0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant s_bottom_right: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant t_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1), 
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1));

constant t_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0));
 








constant t_bottom_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant t_bottom_right: sprite_block :=
((1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),  
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant a_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant a_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),   
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0), 
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0), 
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0));

constant a_bottom_left: sprite_block :=
((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant a_bottom_right: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0), 
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0), 
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant r_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0));

constant r_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0), 
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)); 

constant r_bottom_left: sprite_block :=
((0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant r_bottom_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)); 

constant p_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1));

constant p_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0));

constant p_bottom_left: sprite_block :=
((0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant p_bottom_right: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant e_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant e_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant e_bottom_left: sprite_block :=
((0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant e_bottom_right: sprite_block :=
((1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant c_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0));

constant c_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant c_bottom_left: sprite_block :=
((0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant c_bottom_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant d_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0));

constant d_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0));

constant d_bottom_left: sprite_block :=
((0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant d_bottom_right: sprite_block :=
((0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant exclamation_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1));

constant exclamation_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant exclamation_bottom_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1), 
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1),  
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant exclamation_bottom_right: sprite_block :=
((1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0), 
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));



constant j_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant j_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0));

constant j_bottom_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant j_bottom_right: sprite_block :=
((0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant b_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

constant b_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0));


constant b_bottom_right: sprite_block :=
((1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant b_bottom_left: sprite_block :=
((0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant o_top_right: sprite_block := 
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0));

constant o_top_left: sprite_block := 
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0));


constant o_bottom_right: sprite_block := 
((0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant o_bottom_left: sprite_block := 
((0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant w_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0));

constant w_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1));


constant w_bottom_right: sprite_block :=
((1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant w_bottom_left: sprite_block :=
((0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant n_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0));

constant n_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0));


constant n_bottom_right: sprite_block :=
((0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant n_bottom_left: sprite_block :=
((0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant big_j_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0));

constant big_j_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));



constant big_j_bottom_right: sprite_block :=
((0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant big_j_bottom_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant m_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1));
 
constant m_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0));

constant m_bottom_left: sprite_block :=
((0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1),
(0,0,0,1,1,1,0,0,0,0,0,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant m_bottom_right: sprite_block :=
((1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(1,1,0,0,0,0,1,1,1,1,1,1,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant u_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0));

constant u_top_left: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0));

constant u_bottom_right: sprite_block :=
((0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant u_bottom_left: sprite_block :=
((0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant little_b_top_left: sprite_block :=((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0));

constant little_b_top_right: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0));

constant little_b_bottom_left: sprite_block :=
((0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant little_b_bottom_right: sprite_block :=
((0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


constant slash_top: sprite_block :=
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0));


constant slash_bottom: sprite_block :=
((0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
(0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
(0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0));


constant colon_top: sprite_block := 
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

constant colon_bottom: sprite_block := 
((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

end package sprite_package;
 